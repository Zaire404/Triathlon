// vsrc/include/test_config_pkg.sv
package test_config_pkg;

  import config_pkg::*;

  localparam config_pkg::user_cfg_t TestCfg = '{
      NRET          : unsigned'(4),
      INSTR_PER_FETCH : unsigned'(4),
      XLEN          : unsigned'(32),
      VLEN          : unsigned'(32),
      ILEN          : unsigned'(32),
      BPU_USE_GSHARE : unsigned'(1),
      BPU_USE_TAGE : unsigned'(1),
      BPU_USE_TOURNAMENT : unsigned'(1),
      BPU_BTB_HASH_ENABLE : unsigned'(1),
      BPU_BHT_HASH_ENABLE : unsigned'(1),
      BPU_BTB_ENTRIES : unsigned'(128),
      BPU_BHT_ENTRIES : unsigned'(512),
      BPU_RAS_DEPTH : unsigned'(16),
      BPU_GHR_BITS : unsigned'(8),
      BPU_USE_SC_L : unsigned'(1),
      BPU_SC_L_ENTRIES : unsigned'(1024),
      BPU_SC_L_CONF_THRESH : unsigned'(3),
      BPU_SC_L_REQUIRE_DISAGREE : unsigned'(1),
      BPU_SC_L_REQUIRE_BOTH_WEAK : unsigned'(1),
      BPU_SC_L_BLOCK_ON_TAGE_HIT : unsigned'(0),
      BPU_USE_LOOP : unsigned'(1),
      BPU_LOOP_ENTRIES : unsigned'(128),
      BPU_LOOP_TAG_BITS : unsigned'(10),
      BPU_LOOP_CONF_THRESH : unsigned'(2),
      BPU_USE_ITTAGE : unsigned'(1),
      BPU_ITTAGE_ENTRIES : unsigned'(128),
      BPU_ITTAGE_TAG_BITS : unsigned'(10),
      BPU_TAGE_OVERRIDE_MIN_PROVIDER : unsigned'(2),
      BPU_TAGE_OVERRIDE_REQUIRE_LEGACY_WEAK : unsigned'(1),
      BPU_TAGE_TAG_BITS : unsigned'(8),
      BPU_TAGE_HIST_LEN0 : unsigned'(2),
      BPU_TAGE_HIST_LEN1 : unsigned'(4),
      BPU_TAGE_HIST_LEN2 : unsigned'(8),
      BPU_TAGE_HIST_LEN3 : unsigned'(16),
      BPU_PATH_HIST_BITS : unsigned'(16),
      BPU_TRACK_DEPTH : unsigned'(16),
      ICACHE_HIT_PIPELINE_EN : unsigned'(1),
      IFU_FETCHQ_BYPASS_EN : unsigned'(1),
      IFU_REQ_DEPTH : unsigned'(16),
      IFU_INF_DEPTH : unsigned'(16),
      IFU_FQ_DEPTH : unsigned'(16),
      ENABLE_COMMIT_RAS_UPDATE : unsigned'(1),
      DCACHE_MSHR_SIZE : unsigned'(8),
      RENAME_PENDING_DEPTH : unsigned'(128),
      ROB_DEPTH : unsigned'(128),
      LSU_GROUP_SIZE : unsigned'(4),
      SB_DEPTH : unsigned'(16),
      IBUFFER_DEPTH : unsigned'(16),
      ROB_MAX_COMMIT_BR : unsigned'(1),
      ROB_MAX_COMMIT_ST : unsigned'(1),
      ROB_MAX_COMMIT_LD : unsigned'(2),
      RS_DEPTH     : unsigned'(64),
      ALU_COUNT    : unsigned'(4),
      ICACHE_BYTE_SIZE : unsigned'(8192),
      ICACHE_SET_ASSOC : unsigned'(4),
      ICACHE_LINE_WIDTH : unsigned'(256),

      // DCache (默认与 ICache 同行宽，方便复用 AXI beat 聚合)
      DCACHE_BYTE_SIZE : unsigned'(8192),
      DCACHE_SET_ASSOC : unsigned'(4),
      DCACHE_LINE_WIDTH : unsigned'(256)
  };

endpackage : test_config_pkg
