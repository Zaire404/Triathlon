import config_pkg::*;
import build_config_pkg::*;
import global_config_pkg::*;

module tb_bpu (
    // --- 输入端口  ---
    input logic clk_i,
    input logic rst_i,
    input logic ifu_ready_i,
    input logic ifu_valid_i,
    input logic [Cfg.XLEN - 1:0] pc_i,
    input logic update_valid_i,
    input logic [Cfg.XLEN-1:0] update_pc_i,
    input logic update_is_cond_i,
    input logic update_taken_i,
    input logic [Cfg.XLEN-1:0] update_target_i,
    input logic update_is_call_i,
    input logic update_is_ret_i,
    input logic [Cfg.NRET-1:0] ras_update_valid_i,
    input logic [Cfg.NRET-1:0] ras_update_is_call_i,
    input logic [Cfg.NRET-1:0] ras_update_is_ret_i,
    input logic [Cfg.NRET-1:0][Cfg.PLEN-1:0] ras_update_pc_i,
    input logic flush_i,
    // --- 输出端口  ---
    output logic [Cfg.XLEN-1:0] npc_o,
    output logic pred_slot_valid_o,
    output logic [$clog2(Cfg.INSTR_PER_FETCH)-1:0] pred_slot_idx_o,
    output logic [Cfg.XLEN-1:0] pred_slot_target_o,
    output logic [Cfg.BPU_GHR_BITS-1:0] dbg_ghr_o
);
  // Keep tb_bpu deterministic for legacy hysteresis tests.
  // Frontend integration uses Cfg.BPU_USE_GSHARE.
  localparam bit TB_BPU_USE_GSHARE = 1'b0;
  localparam bit TB_BPU_USE_TAGE = 1'b0;
  localparam bit TB_BPU_USE_ITTAGE = 1'b1;
  localparam int unsigned TB_BPU_BTB_ENTRIES = 128;
  localparam int unsigned TB_BPU_BHT_ENTRIES = 512;
  localparam bit TB_BPU_BTB_HASH_ENABLE = 1'b1;
  localparam bit TB_BPU_BHT_HASH_ENABLE = 1'b1;

  handshake_t  ifu_to_bpu_handshake_i;
  handshake_t  bpu_to_ifu_handshake_o;
  ifu_to_bpu_t ifu_to_bpu_i;
  bpu_to_ifu_t bpu_to_ifu_o;
  assign ifu_to_bpu_i.pc = pc_i;
  assign ifu_to_bpu_handshake_i.ready = ifu_ready_i;
  assign ifu_to_bpu_handshake_i.valid = ifu_valid_i;
  bpu #(
      .Cfg(Cfg),
      .BTB_ENTRIES(TB_BPU_BTB_ENTRIES),
      .BHT_ENTRIES(TB_BPU_BHT_ENTRIES),
      .BTB_HASH_ENABLE(TB_BPU_BTB_HASH_ENABLE),
      .BHT_HASH_ENABLE(TB_BPU_BHT_HASH_ENABLE),
      .USE_GSHARE(TB_BPU_USE_GSHARE),
      .USE_TAGE(TB_BPU_USE_TAGE),
      .USE_ITTAGE(TB_BPU_USE_ITTAGE)
  ) i_BPU (
      .clk_i(clk_i),
      .rst_i(rst_i),
      .ifu_to_bpu_handshake_i(ifu_to_bpu_handshake_i),
      .ifu_to_bpu_i(ifu_to_bpu_i),
      .update_valid_i(update_valid_i),
      .update_pc_i(update_pc_i),
      .update_is_cond_i(update_is_cond_i),
      .update_taken_i(update_taken_i),
      .update_target_i(update_target_i),
      .update_is_call_i(update_is_call_i),
      .update_is_ret_i(update_is_ret_i),
      .ras_update_valid_i(ras_update_valid_i),
      .ras_update_is_call_i(ras_update_is_call_i),
      .ras_update_is_ret_i(ras_update_is_ret_i),
      .ras_update_pc_i(ras_update_pc_i),
      .flush_i(flush_i),

      .bpu_to_ifu_handshake_o(bpu_to_ifu_handshake_o),
      .bpu_to_ifu_o(bpu_to_ifu_o)
  );
  assign npc_o = bpu_to_ifu_o.npc;
  assign pred_slot_valid_o = bpu_to_ifu_o.pred_slot_valid;
  assign pred_slot_idx_o = bpu_to_ifu_o.pred_slot_idx;
  assign pred_slot_target_o = bpu_to_ifu_o.pred_slot_target;
  assign dbg_ghr_o = i_BPU.ghr_q;
endmodule
